-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sun Nov 20 14:33:13 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY maquina_de_estados IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END maquina_de_estados;

ARCHITECTURE BEHAVIOR OF maquina_de_estados IS
    TYPE type_fstate IS (a,b,c,d,e,f,g);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= a;
            Z <= "0000";
        ELSE
            Z <= "0000";
            CASE fstate IS
                WHEN a =>
                    IF ((x = '0')) THEN
                        reg_fstate <= b;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= e;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= a;
                    END IF;

                    Z <= "0000";
                WHEN b =>
                    reg_fstate <= c;

                    Z <= "0110";
                WHEN c =>
                    IF ((x = '0')) THEN
                        reg_fstate <= d;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= g;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= c;
                    END IF;

                    Z <= "1111";
                WHEN d =>
                    reg_fstate <= a;

                    Z <= "1001";
                WHEN e =>
                    reg_fstate <= f;

                    Z <= "1000";
                WHEN f =>
                    reg_fstate <= g;

                    Z <= "1100";
                WHEN g =>
                    reg_fstate <= a;

                    Z <= "1110";
                WHEN OTHERS => 
                    Z <= "XXXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
