library verilog;
use verilog.vl_types.all;
entity maquina_de_estados_vlg_vec_tst is
end maquina_de_estados_vlg_vec_tst;
