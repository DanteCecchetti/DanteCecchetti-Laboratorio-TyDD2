library verilog;
use verilog.vl_types.all;
entity ParteDb_vlg_vec_tst is
end ParteDb_vlg_vec_tst;
