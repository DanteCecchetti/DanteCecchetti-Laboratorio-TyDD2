library verilog;
use verilog.vl_types.all;
entity Sum4bit_vlg_vec_tst is
end Sum4bit_vlg_vec_tst;
