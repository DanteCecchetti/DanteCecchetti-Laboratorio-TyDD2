library verilog;
use verilog.vl_types.all;
entity sumador_FFD_vlg_vec_tst is
end sumador_FFD_vlg_vec_tst;
